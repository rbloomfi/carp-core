`ifndef MEMORY_LAYOUT_SVH
`define MEMORY_LAYOUT_SVH

parameter DATA_BASE_ADDR = 14'h6000;
`endif

