`timescale 1ns/1ps

module tb_MUL();

    logic [31:0] RS1_E, RS1_M, RS1_W;
    logic [31:0] RS2_E, RS2_M, RS2_W;

    typedef struct packed {
        logic SIGN,
        logic CYCLES,
        logic OP,
          
    } struct_name;

endmodule